bind BranchCondition_clk checker_branch chk_branch(.*);