bind BranchCondition checker_branch chk_branch(.*);