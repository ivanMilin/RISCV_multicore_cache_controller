bind ImmediateGenerator checker_imm_gen chk_imm_gen(.*);