bind top ref_model_top chk_ref_model_top(.*);
