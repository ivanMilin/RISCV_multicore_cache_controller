bind Top ref_model_top chk_ref_model_top(.*);
