bind Controller checker_controller chk_controller(.*);
