bind Processor ref_model chk_ref_model(.*);
