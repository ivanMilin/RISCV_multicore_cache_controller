`define TYPE_R 7'b0110011
`define TYPE_I 7'b0010011
`define TYPE_L 7'b0000011
`define TYPE_S 7'b0100011
`define TYPE_B 7'b1100011
`define TYPE_U 7'b0110111
`define TYPE_J 7'b1101111
